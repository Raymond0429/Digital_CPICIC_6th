module matrix_cal_top 
#(parameter DATA_WIDTH = 'd128)
(   input clk         ,
    input rst_n       ,
    input src_row_vld ,
    input src_row_rdy ,
    input [DATA_WIDTH*16-1:0] src_row_data,

    output tmp_col_vld ,
    output tmp_col_rdy ,
    output [(DATA_WIDTH+4)*16-1:0] tmp_col_data
 );




endmodule